----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 03/31/2021 07:24:23 PM
-- Design Name: 
-- Module Name: top - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;
use ieee.std_logic_unsigned.all;
use IEEE.math_real.all;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

library xil_defaultlib;
use xil_defaultlib.math_functions.all;
use xil_defaultlib.firmware_config.all;
use xil_defaultlib.packet_defs.all;
use xil_defaultlib.fox_defs.all;

entity board_top is
    Port ( 
           CPU_RESETN   : in STD_LOGIC;
           clk          : in STD_LOGIC;
           LED          : out STD_LOGIC_VECTOR(3 downto 0);
           UART_RXD_OUT : out std_logic
    );
end board_top;

architecture Behavioral of board_top is

    component top
        generic (
            -- Fox's algorithm network paramters
            FOX_NETWORK_STAGES  : integer := 2;
            FOX_NETWORK_NODES   : integer := 4;
            
            FOX_FIRMWARE            : string := "firmware_hoplite.hex";
            FOX_FIRMWARE_MEM_SIZE   : integer := 4096; 
            
            RESULT_FIRMWARE             : string := "firmware_hoplite_result.hex";
            RESULT_FIRMWARE_MEM_SIZE    : integer := 8192;
            
            CLK_FREQ            : integer := 50e6;
            ENABLE_UART         : boolean := False
        );
        port (
            clk                 : in std_logic;
            reset_n             : in std_logic;
            
            LED                 : out STD_LOGIC_VECTOR((FOX_NETWORK_NODES-1) downto 0);
            
            out_char            : out t_Char;
            out_char_en         : out t_MessageValid;
            
            uart_tx             : out std_logic;
            
            out_matrix          : out t_MatrixOut;
            out_matrix_en       : out t_MessageValid;
            out_matrix_end_row  : out t_MessageValid;
            out_matrix_end      : out t_MessageValid;
            
            ila_multicast_out        : out std_logic_vector((BUS_WIDTH-1) downto 0);
            ila_multicast_out_valid  : out std_logic;
            
            ila_x_out            : out std_logic_vector((BUS_WIDTH-1) downto 0);
            ila_x_out_valid      : out std_logic;
           
            ila_y_out            : out std_logic_vector((BUS_WIDTH-1) downto 0);
            ila_y_out_valid      : out std_logic
        );
    end component top;
    
    component clock_divider 
        Port ( 
            CLK_50MHZ   : out STD_LOGIC;
            reset       : in STD_LOGIC;
            locked      : out STD_LOGIC;
            clk_in1     : in STD_LOGIC
        );
    end component clock_divider;
        
    signal reset    : std_logic;
    signal locked   : std_logic;
        
    signal clkdiv2  : std_logic;
        
    constant CLK_FREQ       : integer := 50e6;
    constant ENABLE_UART    : boolean := True;
    
    signal reset_n  : std_logic;

    component multicast_ila
        Port (
            clk : in std_logic;
           
            probe0  : in std_logic_vector(58 downto 0);
            probe1  : in std_logic_vector(0 downto 0)
        );
    end component multicast_ila;
    
    constant ENABLE_MULTICAST_ROUTER_0_ILA : boolean := True;
    
    signal ila_multicast_out        : std_logic_vector((BUS_WIDTH-1) downto 0);
    signal ila_multicast_out_valid  : std_logic;
    
    component hoplite_router_ila
        Port (
            clk : in std_logic;
           
            probe0  : in std_logic_vector(58 downto 0);
            probe1  : in std_logic_vector(0 downto 0);
            
            probe2  : in std_logic_vector(58 downto 0);
            probe3  : in std_logic_vector(0 downto 0)
        );
    end component hoplite_router_ila;
    
    constant ENABLE_HOPLITE_ROUTER_0_ILA : boolean := True;
    
    signal ila_x_out        : std_logic_vector((BUS_WIDTH-1) downto 0);
    signal ila_x_out_valid  : std_logic;
    
    signal ila_y_out        : std_logic_vector((BUS_WIDTH-1) downto 0);
    signal ila_y_out_valid  : std_logic;

begin

    reset   <= not CPU_RESETN;

    -- Clock divider
    DIVIDER: clock_divider
        port map (
            clk_in1     => clk,
            reset       => reset,
            locked      => locked,
            CLK_50MHZ   => clkdiv2
        );
    
    reset_n <= CPU_RESETN and locked;

    FOX_TOP: top
        generic map (
            FOX_NETWORK_STAGES  => FOX_NETWORK_STAGES,
            FOX_NETWORK_NODES   => FOX_NETWORK_NODES,
            
            FOX_FIRMWARE            => FOX_FIRMWARE,
            FOX_FIRMWARE_MEM_SIZE   => FOX_MEM_SIZE,
            
            RESULT_FIRMWARE             => RESULT_FIRMWARE,
            RESULT_FIRMWARE_MEM_SIZE    => RESULT_MEM_SIZE,
            
            CLK_FREQ            => CLK_FREQ,
            ENABLE_UART         => ENABLE_UART
        )
        port map (
            clk                 => clkdiv2,
            reset_n             => reset_n,
            
            LED                 => LED,
            
            out_char            => open,
            out_char_en         => open,
            
            uart_tx             => UART_RXD_OUT,
            
            out_matrix          => open,
            out_matrix_en       => open,
            out_matrix_end_row  => open,
            out_matrix_end      => open,
            
            ila_multicast_out       => ila_multicast_out,
            ila_multicast_out_valid => ila_multicast_out_valid,
            
            ila_x_out           => ila_x_out,
            ila_x_out_valid     => ila_x_out_valid,
            
            ila_y_out           => ila_y_out,
            ila_y_out_valid     => ila_y_out_valid
        );
      
    MULTICAST_ROUTER_0_ILA_GEN: if (ENABLE_MULTICAST_ROUTER_0_ILA = True) generate  
        MULTICAST_ROUTER_0_ILA: multicast_ila
            port map (
                clk         => clkdiv2,
               
                probe0      => ila_multicast_out,
                probe1(0)   => ila_multicast_out_valid
            );
    end generate MULTICAST_ROUTER_0_ILA_GEN;
    
    HOPLITE_ROUTER_0_ILA_GEN: if (ENABLE_HOPLITE_ROUTER_0_ILA = True) generate  
        HOPLITE_ROUTER_0_ILA: hoplite_router_ila
            port map (
                clk         => clkdiv2,
               
                probe0      => ila_x_out,
                probe1(0)   => ila_x_out_valid,
                
                probe2      => ila_y_out,
                probe3(0)   => ila_y_out_valid
            );
    end generate HOPLITE_ROUTER_0_ILA_GEN;

end Behavioral;
