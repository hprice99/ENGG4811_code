`ifndef IO_VH
`define IO_VH

// Character output
`define CHAR_OUTPUT      32'h1000_0000
`define CHAR_OUTPUT_READY_INPUT      32'h1000_0010




// Node details
`define MATRIX_INIT_FROM_FILE_INPUT      32'h5000_0000

// Matrix
`define MATRIX_OUTPUT      32'h6000_0000
`define MATRIX_END_ROW_OUTPUT      32'h6000_0010
`define MATRIX_END_OUTPUT      32'h6000_0020
`define MATRIX_INIT_TYPE_INPUT      32'h6000_0030
`define MATRIX_INIT_X_COORD_INPUT      32'h6000_0040
`define MATRIX_INIT_Y_COORD_INPUT      32'h6000_0050
`define MATRIX_INIT_ELEMENT_INPUT      32'h6000_0060
`define MATRIX_INIT_READ_OUTPUT      32'h6000_0070
`define MATRIX_MULTIPLY_DONE_OUTPUT      32'h6000_0080


`endif