library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

package firmware_config is 

    constant FOX_FIRMWARE       : string := "firmware_fox_hoplite_multicast.hex";
    constant FOX_MEM_SIZE       : integer := 4096;

    constant RESULT_FIRMWARE    : string := "firmware_fox_hoplite_multicast_result.hex";
    constant RESULT_MEM_SIZE    : integer := 8192;

end package firmware_config;

package body firmware_config is

end package body firmware_config;