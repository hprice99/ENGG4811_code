library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

package firmware_config is 

    constant FOX_FIRMWARE       : string := "firmware_single_core.hex";
    constant FOX_MEM_SIZE       : integer := 32678;


end package firmware_config;

package body firmware_config is

end package body firmware_config;